-------------------------------------------------------------------------------
-- Title      : sigmoid
-- Project    : SNN
-------------------------------------------------------------------------------
-- File       : sigmoid.vhd
-- Author     : Isadora Sophia e Matheus Diamantino
-- Company    : Unicamp!
-- Created    : 2016-06-11
-- Last update: 2016-06-11
-- Platform   : Cyclone II
-- Standard   : VHDL'2008
-------------------------------------------------------------------------------
-- Description: Sigmoid function, implemented with a lookup table
-------------------------------------------------------------------------------
-- Copyright (c) 2016
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  							Description
-- 2016-06-11  0.1      Isadora Sophia e Matheus Diamantino	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- fixed point lib
library work;
use work.fixed_pkg.all;

-- our own lib
use work.extra_pkg.all;

entity sigmoid is
    port (
		i: in  sfixed(dec - 1 downto -frac);
		o: out sfixed(dec - 1 downto -frac)
	);
end sigmoid;

architecture lut of sigmoid is
	subtype temp is std_logic_vector(i'length - 1 downto 0); -- in order to convert sfixed to std_logic_vector
	signal t_i, t_o : temp;
begin
	-- convert input to std_logic
	t_i <= temp(i);
	
	-- convert output back to sfixed
	o <= to_sfixed(t_o, o'high, o'low);
	
	-- lookup table
	t_o <=
		"0000000100000000" when to_integer(signed(t_i(i'length - 1 downto 3))) > 553 else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0001000000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111110000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000111000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110110000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000110000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101110000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000101000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100110000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000100000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011110000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011101000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011100000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011011000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011010000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011001000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000011000000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111001" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010111000" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110111" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110110" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110101" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110100" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110011" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110010" else
		"0000000011111111" when t_i(i'length - 1 downto 3) = "0000010110001" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010110000" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101111" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101110" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101101" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101100" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101011" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101010" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101001" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010101000" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100111" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100110" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100101" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100100" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100011" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100010" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100001" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010100000" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010011111" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010011110" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010011101" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010011100" else
		"0000000011111110" when t_i(i'length - 1 downto 3) = "0000010011011" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010011010" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010011001" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010011000" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010111" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010110" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010101" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010100" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010011" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010010" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010001" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010010000" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010001111" else
		"0000000011111101" when t_i(i'length - 1 downto 3) = "0000010001110" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001101" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001100" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001011" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001010" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001001" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010001000" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010000111" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010000110" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010000101" else
		"0000000011111100" when t_i(i'length - 1 downto 3) = "0000010000100" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000010000011" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000010000010" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000010000001" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000010000000" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000001111111" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000001111110" else
		"0000000011111011" when t_i(i'length - 1 downto 3) = "0000001111101" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001111100" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001111011" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001111010" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001111001" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001111000" else
		"0000000011111010" when t_i(i'length - 1 downto 3) = "0000001110111" else
		"0000000011111001" when t_i(i'length - 1 downto 3) = "0000001110110" else
		"0000000011111001" when t_i(i'length - 1 downto 3) = "0000001110101" else
		"0000000011111001" when t_i(i'length - 1 downto 3) = "0000001110100" else
		"0000000011111001" when t_i(i'length - 1 downto 3) = "0000001110011" else
		"0000000011111001" when t_i(i'length - 1 downto 3) = "0000001110010" else
		"0000000011111000" when t_i(i'length - 1 downto 3) = "0000001110001" else
		"0000000011111000" when t_i(i'length - 1 downto 3) = "0000001110000" else
		"0000000011111000" when t_i(i'length - 1 downto 3) = "0000001101111" else
		"0000000011111000" when t_i(i'length - 1 downto 3) = "0000001101110" else
		"0000000011110111" when t_i(i'length - 1 downto 3) = "0000001101101" else
		"0000000011110111" when t_i(i'length - 1 downto 3) = "0000001101100" else
		"0000000011110111" when t_i(i'length - 1 downto 3) = "0000001101011" else
		"0000000011110111" when t_i(i'length - 1 downto 3) = "0000001101010" else
		"0000000011110110" when t_i(i'length - 1 downto 3) = "0000001101001" else
		"0000000011110110" when t_i(i'length - 1 downto 3) = "0000001101000" else
		"0000000011110110" when t_i(i'length - 1 downto 3) = "0000001100111" else
		"0000000011110110" when t_i(i'length - 1 downto 3) = "0000001100110" else
		"0000000011110101" when t_i(i'length - 1 downto 3) = "0000001100101" else
		"0000000011110101" when t_i(i'length - 1 downto 3) = "0000001100100" else
		"0000000011110101" when t_i(i'length - 1 downto 3) = "0000001100011" else
		"0000000011110100" when t_i(i'length - 1 downto 3) = "0000001100010" else
		"0000000011110100" when t_i(i'length - 1 downto 3) = "0000001100001" else
		"0000000011110100" when t_i(i'length - 1 downto 3) = "0000001100000" else
		"0000000011110011" when t_i(i'length - 1 downto 3) = "0000001011111" else
		"0000000011110011" when t_i(i'length - 1 downto 3) = "0000001011110" else
		"0000000011110011" when t_i(i'length - 1 downto 3) = "0000001011101" else
		"0000000011110010" when t_i(i'length - 1 downto 3) = "0000001011100" else
		"0000000011110010" when t_i(i'length - 1 downto 3) = "0000001011011" else
		"0000000011110001" when t_i(i'length - 1 downto 3) = "0000001011010" else
		"0000000011110001" when t_i(i'length - 1 downto 3) = "0000001011001" else
		"0000000011110001" when t_i(i'length - 1 downto 3) = "0000001011000" else
		"0000000011110000" when t_i(i'length - 1 downto 3) = "0000001010111" else
		"0000000011110000" when t_i(i'length - 1 downto 3) = "0000001010110" else
		"0000000011101111" when t_i(i'length - 1 downto 3) = "0000001010101" else
		"0000000011101111" when t_i(i'length - 1 downto 3) = "0000001010100" else
		"0000000011101110" when t_i(i'length - 1 downto 3) = "0000001010011" else
		"0000000011101110" when t_i(i'length - 1 downto 3) = "0000001010010" else
		"0000000011101101" when t_i(i'length - 1 downto 3) = "0000001010001" else
		"0000000011101101" when t_i(i'length - 1 downto 3) = "0000001010000" else
		"0000000011101100" when t_i(i'length - 1 downto 3) = "0000001001111" else
		"0000000011101011" when t_i(i'length - 1 downto 3) = "0000001001110" else
		"0000000011101011" when t_i(i'length - 1 downto 3) = "0000001001101" else
		"0000000011101010" when t_i(i'length - 1 downto 3) = "0000001001100" else
		"0000000011101010" when t_i(i'length - 1 downto 3) = "0000001001011" else
		"0000000011101001" when t_i(i'length - 1 downto 3) = "0000001001010" else
		"0000000011101000" when t_i(i'length - 1 downto 3) = "0000001001001" else
		"0000000011101000" when t_i(i'length - 1 downto 3) = "0000001001000" else
		"0000000011100111" when t_i(i'length - 1 downto 3) = "0000001000111" else
		"0000000011100110" when t_i(i'length - 1 downto 3) = "0000001000110" else
		"0000000011100110" when t_i(i'length - 1 downto 3) = "0000001000101" else
		"0000000011100101" when t_i(i'length - 1 downto 3) = "0000001000100" else
		"0000000011100100" when t_i(i'length - 1 downto 3) = "0000001000011" else
		"0000000011100011" when t_i(i'length - 1 downto 3) = "0000001000010" else
		"0000000011100011" when t_i(i'length - 1 downto 3) = "0000001000001" else
		"0000000011100010" when t_i(i'length - 1 downto 3) = "0000001000000" else
		"0000000011100001" when t_i(i'length - 1 downto 3) = "0000000111111" else
		"0000000011100000" when t_i(i'length - 1 downto 3) = "0000000111110" else
		"0000000011011111" when t_i(i'length - 1 downto 3) = "0000000111101" else
		"0000000011011110" when t_i(i'length - 1 downto 3) = "0000000111100" else
		"0000000011011101" when t_i(i'length - 1 downto 3) = "0000000111011" else
		"0000000011011100" when t_i(i'length - 1 downto 3) = "0000000111010" else
		"0000000011011011" when t_i(i'length - 1 downto 3) = "0000000111001" else
		"0000000011011010" when t_i(i'length - 1 downto 3) = "0000000111000" else
		"0000000011011001" when t_i(i'length - 1 downto 3) = "0000000110111" else
		"0000000011011000" when t_i(i'length - 1 downto 3) = "0000000110110" else
		"0000000011010111" when t_i(i'length - 1 downto 3) = "0000000110101" else
		"0000000011010110" when t_i(i'length - 1 downto 3) = "0000000110100" else
		"0000000011010101" when t_i(i'length - 1 downto 3) = "0000000110011" else
		"0000000011010100" when t_i(i'length - 1 downto 3) = "0000000110010" else
		"0000000011010011" when t_i(i'length - 1 downto 3) = "0000000110001" else
		"0000000011010010" when t_i(i'length - 1 downto 3) = "0000000110000" else
		"0000000011010001" when t_i(i'length - 1 downto 3) = "0000000101111" else
		"0000000011001111" when t_i(i'length - 1 downto 3) = "0000000101110" else
		"0000000011001110" when t_i(i'length - 1 downto 3) = "0000000101101" else
		"0000000011001101" when t_i(i'length - 1 downto 3) = "0000000101100" else
		"0000000011001100" when t_i(i'length - 1 downto 3) = "0000000101011" else
		"0000000011001010" when t_i(i'length - 1 downto 3) = "0000000101010" else
		"0000000011001001" when t_i(i'length - 1 downto 3) = "0000000101001" else
		"0000000011001000" when t_i(i'length - 1 downto 3) = "0000000101000" else
		"0000000011000110" when t_i(i'length - 1 downto 3) = "0000000100111" else
		"0000000011000101" when t_i(i'length - 1 downto 3) = "0000000100110" else
		"0000000011000011" when t_i(i'length - 1 downto 3) = "0000000100101" else
		"0000000011000010" when t_i(i'length - 1 downto 3) = "0000000100100" else
		"0000000011000001" when t_i(i'length - 1 downto 3) = "0000000100011" else
		"0000000010111111" when t_i(i'length - 1 downto 3) = "0000000100010" else
		"0000000010111110" when t_i(i'length - 1 downto 3) = "0000000100001" else
		"0000000010111100" when t_i(i'length - 1 downto 3) = "0000000100000" else
		"0000000010111010" when t_i(i'length - 1 downto 3) = "0000000011111" else
		"0000000010111001" when t_i(i'length - 1 downto 3) = "0000000011110" else
		"0000000010110111" when t_i(i'length - 1 downto 3) = "0000000011101" else
		"0000000010110110" when t_i(i'length - 1 downto 3) = "0000000011100" else
		"0000000010110100" when t_i(i'length - 1 downto 3) = "0000000011011" else
		"0000000010110010" when t_i(i'length - 1 downto 3) = "0000000011010" else
		"0000000010110001" when t_i(i'length - 1 downto 3) = "0000000011001" else
		"0000000010101111" when t_i(i'length - 1 downto 3) = "0000000011000" else
		"0000000010101101" when t_i(i'length - 1 downto 3) = "0000000010111" else
		"0000000010101011" when t_i(i'length - 1 downto 3) = "0000000010110" else
		"0000000010101010" when t_i(i'length - 1 downto 3) = "0000000010101" else
		"0000000010101000" when t_i(i'length - 1 downto 3) = "0000000010100" else
		"0000000010100110" when t_i(i'length - 1 downto 3) = "0000000010011" else
		"0000000010100100" when t_i(i'length - 1 downto 3) = "0000000010010" else
		"0000000010100010" when t_i(i'length - 1 downto 3) = "0000000010001" else
		"0000000010100000" when t_i(i'length - 1 downto 3) = "0000000010000" else
		"0000000010011111" when t_i(i'length - 1 downto 3) = "0000000001111" else
		"0000000010011101" when t_i(i'length - 1 downto 3) = "0000000001110" else
		"0000000010011011" when t_i(i'length - 1 downto 3) = "0000000001101" else
		"0000000010011001" when t_i(i'length - 1 downto 3) = "0000000001100" else
		"0000000010010111" when t_i(i'length - 1 downto 3) = "0000000001011" else
		"0000000010010101" when t_i(i'length - 1 downto 3) = "0000000001010" else
		"0000000010010011" when t_i(i'length - 1 downto 3) = "0000000001001" else
		"0000000010010001" when t_i(i'length - 1 downto 3) = "0000000001000" else
		"0000000010001111" when t_i(i'length - 1 downto 3) = "0000000000111" else
		"0000000010001101" when t_i(i'length - 1 downto 3) = "0000000000110" else
		"0000000010001011" when t_i(i'length - 1 downto 3) = "0000000000101" else
		"0000000010001001" when t_i(i'length - 1 downto 3) = "0000000000100" else
		"0000000010000111" when t_i(i'length - 1 downto 3) = "0000000000011" else
		"0000000010000101" when t_i(i'length - 1 downto 3) = "0000000000010" else
		"0000000010000011" when t_i(i'length - 1 downto 3) = "0000000000001" else
		"0000000010000001" when t_i(i'length - 1 downto 3) = "0000000000000" else
		"0000000001111111" when t_i(i'length - 1 downto 3) = "1111111111111" else
		"0000000001111101" when t_i(i'length - 1 downto 3) = "1000000000000" else
		"0000000001111011" when t_i(i'length - 1 downto 3) = "1000000000001" else
		"0000000001111001" when t_i(i'length - 1 downto 3) = "1000000000010" else
		"0000000001110111" when t_i(i'length - 1 downto 3) = "1000000000011" else
		"0000000001110101" when t_i(i'length - 1 downto 3) = "1000000000100" else
		"0000000001110011" when t_i(i'length - 1 downto 3) = "1000000000101" else
		"0000000001110001" when t_i(i'length - 1 downto 3) = "1000000000110" else
		"0000000001101111" when t_i(i'length - 1 downto 3) = "1000000000111" else
		"0000000001101101" when t_i(i'length - 1 downto 3) = "1000000001000" else
		"0000000001101011" when t_i(i'length - 1 downto 3) = "1000000001001" else
		"0000000001101001" when t_i(i'length - 1 downto 3) = "1000000001010" else
		"0000000001101000" when t_i(i'length - 1 downto 3) = "1000000001011" else
		"0000000001100110" when t_i(i'length - 1 downto 3) = "1000000001100" else
		"0000000001100100" when t_i(i'length - 1 downto 3) = "1000000001101" else
		"0000000001100010" when t_i(i'length - 1 downto 3) = "1000000001110" else
		"0000000001100000" when t_i(i'length - 1 downto 3) = "1000000001111" else
		"0000000001011110" when t_i(i'length - 1 downto 3) = "1000000010000" else
		"0000000001011100" when t_i(i'length - 1 downto 3) = "1000000010001" else
		"0000000001011010" when t_i(i'length - 1 downto 3) = "1000000010010" else
		"0000000001011001" when t_i(i'length - 1 downto 3) = "1000000010011" else
		"0000000001010111" when t_i(i'length - 1 downto 3) = "1000000010100" else
		"0000000001010101" when t_i(i'length - 1 downto 3) = "1000000010101" else
		"0000000001010011" when t_i(i'length - 1 downto 3) = "1000000010110" else
		"0000000001010001" when t_i(i'length - 1 downto 3) = "1000000010111" else
		"0000000001010000" when t_i(i'length - 1 downto 3) = "1000000011000" else
		"0000000001001110" when t_i(i'length - 1 downto 3) = "1000000011001" else
		"0000000001001100" when t_i(i'length - 1 downto 3) = "1000000011010" else
		"0000000001001011" when t_i(i'length - 1 downto 3) = "1000000011011" else
		"0000000001001001" when t_i(i'length - 1 downto 3) = "1000000011100" else
		"0000000001000111" when t_i(i'length - 1 downto 3) = "1000000011101" else
		"0000000001000110" when t_i(i'length - 1 downto 3) = "1000000011110" else
		"0000000001000100" when t_i(i'length - 1 downto 3) = "1000000011111" else
		"0000000001000011" when t_i(i'length - 1 downto 3) = "1000000100000" else
		"0000000001000001" when t_i(i'length - 1 downto 3) = "1000000100001" else
		"0000000001000000" when t_i(i'length - 1 downto 3) = "1000000100010" else
		"0000000000111110" when t_i(i'length - 1 downto 3) = "1000000100011" else
		"0000000000111101" when t_i(i'length - 1 downto 3) = "1000000100100" else
		"0000000000111011" when t_i(i'length - 1 downto 3) = "1000000100101" else
		"0000000000111010" when t_i(i'length - 1 downto 3) = "1000000100110" else
		"0000000000111000" when t_i(i'length - 1 downto 3) = "1000000100111" else
		"0000000000110111" when t_i(i'length - 1 downto 3) = "1000000101000" else
		"0000000000110110" when t_i(i'length - 1 downto 3) = "1000000101001" else
		"0000000000110100" when t_i(i'length - 1 downto 3) = "1000000101010" else
		"0000000000110011" when t_i(i'length - 1 downto 3) = "1000000101011" else
		"0000000000110010" when t_i(i'length - 1 downto 3) = "1000000101100" else
		"0000000000110000" when t_i(i'length - 1 downto 3) = "1000000101101" else
		"0000000000101111" when t_i(i'length - 1 downto 3) = "1000000101110" else
		"0000000000101110" when t_i(i'length - 1 downto 3) = "1000000101111" else
		"0000000000101101" when t_i(i'length - 1 downto 3) = "1000000110000" else
		"0000000000101100" when t_i(i'length - 1 downto 3) = "1000000110001" else
		"0000000000101011" when t_i(i'length - 1 downto 3) = "1000000110010" else
		"0000000000101001" when t_i(i'length - 1 downto 3) = "1000000110011" else
		"0000000000101000" when t_i(i'length - 1 downto 3) = "1000000110100" else
		"0000000000100111" when t_i(i'length - 1 downto 3) = "1000000110101" else
		"0000000000100110" when t_i(i'length - 1 downto 3) = "1000000110110" else
		"0000000000100101" when t_i(i'length - 1 downto 3) = "1000000110111" else
		"0000000000100100" when t_i(i'length - 1 downto 3) = "1000000111000" else
		"0000000000100011" when t_i(i'length - 1 downto 3) = "1000000111001" else
		"0000000000100010" when t_i(i'length - 1 downto 3) = "1000000111010" else
		"0000000000100001" when t_i(i'length - 1 downto 3) = "1000000111011" else
		"0000000000100001" when t_i(i'length - 1 downto 3) = "1000000111100" else
		"0000000000100000" when t_i(i'length - 1 downto 3) = "1000000111101" else
		"0000000000011111" when t_i(i'length - 1 downto 3) = "1000000111110" else
		"0000000000011110" when t_i(i'length - 1 downto 3) = "1000000111111" else
		"0000000000011101" when t_i(i'length - 1 downto 3) = "1000001000000" else
		"0000000000011100" when t_i(i'length - 1 downto 3) = "1000001000001" else
		"0000000000011011" when t_i(i'length - 1 downto 3) = "1000001000010" else
		"0000000000011011" when t_i(i'length - 1 downto 3) = "1000001000011" else
		"0000000000011010" when t_i(i'length - 1 downto 3) = "1000001000100" else
		"0000000000011001" when t_i(i'length - 1 downto 3) = "1000001000101" else
		"0000000000011001" when t_i(i'length - 1 downto 3) = "1000001000110" else
		"0000000000011000" when t_i(i'length - 1 downto 3) = "1000001000111" else
		"0000000000010111" when t_i(i'length - 1 downto 3) = "1000001001000" else
		"0000000000010110" when t_i(i'length - 1 downto 3) = "1000001001001" else
		"0000000000010110" when t_i(i'length - 1 downto 3) = "1000001001010" else
		"0000000000010101" when t_i(i'length - 1 downto 3) = "1000001001011" else
		"0000000000010101" when t_i(i'length - 1 downto 3) = "1000001001100" else
		"0000000000010100" when t_i(i'length - 1 downto 3) = "1000001001101" else
		"0000000000010011" when t_i(i'length - 1 downto 3) = "1000001001110" else
		"0000000000010011" when t_i(i'length - 1 downto 3) = "1000001001111" else
		"0000000000010010" when t_i(i'length - 1 downto 3) = "1000001010000" else
		"0000000000010010" when t_i(i'length - 1 downto 3) = "1000001010001" else
		"0000000000010001" when t_i(i'length - 1 downto 3) = "1000001010010" else
		"0000000000010001" when t_i(i'length - 1 downto 3) = "1000001010011" else
		"0000000000010000" when t_i(i'length - 1 downto 3) = "1000001010100" else
		"0000000000010000" when t_i(i'length - 1 downto 3) = "1000001010101" else
		"0000000000001111" when t_i(i'length - 1 downto 3) = "1000001010110" else
		"0000000000001111" when t_i(i'length - 1 downto 3) = "1000001010111" else
		"0000000000001110" when t_i(i'length - 1 downto 3) = "1000001011000" else
		"0000000000001110" when t_i(i'length - 1 downto 3) = "1000001011001" else
		"0000000000001110" when t_i(i'length - 1 downto 3) = "1000001011010" else
		"0000000000001101" when t_i(i'length - 1 downto 3) = "1000001011011" else
		"0000000000001101" when t_i(i'length - 1 downto 3) = "1000001011100" else
		"0000000000001100" when t_i(i'length - 1 downto 3) = "1000001011101" else
		"0000000000001100" when t_i(i'length - 1 downto 3) = "1000001011110" else
		"0000000000001100" when t_i(i'length - 1 downto 3) = "1000001011111" else
		"0000000000001011" when t_i(i'length - 1 downto 3) = "1000001100000" else
		"0000000000001011" when t_i(i'length - 1 downto 3) = "1000001100001" else
		"0000000000001011" when t_i(i'length - 1 downto 3) = "1000001100010" else
		"0000000000001010" when t_i(i'length - 1 downto 3) = "1000001100011" else
		"0000000000001010" when t_i(i'length - 1 downto 3) = "1000001100100" else
		"0000000000001010" when t_i(i'length - 1 downto 3) = "1000001100101" else
		"0000000000001001" when t_i(i'length - 1 downto 3) = "1000001100110" else
		"0000000000001001" when t_i(i'length - 1 downto 3) = "1000001100111" else
		"0000000000001001" when t_i(i'length - 1 downto 3) = "1000001101000" else
		"0000000000001000" when t_i(i'length - 1 downto 3) = "1000001101001" else
		"0000000000001000" when t_i(i'length - 1 downto 3) = "1000001101010" else
		"0000000000001000" when t_i(i'length - 1 downto 3) = "1000001101011" else
		"0000000000001000" when t_i(i'length - 1 downto 3) = "1000001101100" else
		"0000000000000111" when t_i(i'length - 1 downto 3) = "1000001101101" else
		"0000000000000111" when t_i(i'length - 1 downto 3) = "1000001101110" else
		"0000000000000111" when t_i(i'length - 1 downto 3) = "1000001101111" else
		"0000000000000111" when t_i(i'length - 1 downto 3) = "1000001110000" else
		"0000000000000111" when t_i(i'length - 1 downto 3) = "1000001110001" else
		"0000000000000110" when t_i(i'length - 1 downto 3) = "1000001110010" else
		"0000000000000110" when t_i(i'length - 1 downto 3) = "1000001110011" else
		"0000000000000110" when t_i(i'length - 1 downto 3) = "1000001110100" else
		"0000000000000110" when t_i(i'length - 1 downto 3) = "1000001110101" else
		"0000000000000110" when t_i(i'length - 1 downto 3) = "1000001110110" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001110111" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001111000" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001111001" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001111010" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001111011" else
		"0000000000000101" when t_i(i'length - 1 downto 3) = "1000001111100" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000001111101" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000001111110" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000001111111" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000010000000" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000010000001" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000010000010" else
		"0000000000000100" when t_i(i'length - 1 downto 3) = "1000010000011" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010000100" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010000101" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010000110" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010000111" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010001000" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010001001" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010001010" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010001011" else
		"0000000000000011" when t_i(i'length - 1 downto 3) = "1000010001100" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010001101" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010001110" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010001111" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010000" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010001" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010010" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010011" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010100" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010101" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010110" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010010111" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010011000" else
		"0000000000000010" when t_i(i'length - 1 downto 3) = "1000010011001" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011010" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011011" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011100" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011101" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011110" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010011111" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100000" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100001" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100010" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100011" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100100" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100101" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100110" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010100111" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101000" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101001" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101010" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101011" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101100" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101101" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101110" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010101111" else
		"0000000000000001" when t_i(i'length - 1 downto 3) = "1000010110000" else
		"0000000000000000";

end lut;
